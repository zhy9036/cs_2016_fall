

module sram
(
//DE1 board interface
input  wire clk ,
input  wire [2:0] key ,  //buttons = write, read, reset_n
output wire [7:0] ledr,
output wire [7:0] ledg,

// sram signals
output wire [17:0] sram_addr ,
output wire sram_oe_n, sram_we_n,
inout  wire [15:0] sram_dq,
output wire sram_ce_n , sram_lb_n, sram_ub_n
);


//internal signals
reg [2:0] state_reg, state_next;
reg [17:0] count_reg, count_next;
wire  reset_n = key[0];
wire  read  = key[1];
wire  write = key[2];
reg   start_n;
reg   rw;
wire ready ;
wire [15:0] data_read;
wire pulse;
reg rst_pulse;

localparam [2:0] state_idle    = 3'b000, // states
						state_read1  = 3'b001,
						state_read2  = 3'b010,
						state_write1 = 3'b011,
						state_write2 = 3'b100;
//SRAM CONTROLLER
sram_ctrl device0(.clk(clk), .reset_n(reset_n), .start_n(start_n), .rw(rw), .addr_in(count_reg), .data_write(count_reg[15:0]), .ready(ready),
					.data_read(data_read), .sram_addr(sram_addr), .we_n(sram_we_n), .oe_n(sram_oe_n), 
					.data_io(sram_dq), .ce_a_n(sram_ce_n), .ub_a_n(sram_ub_n), .lb_a_n(sram_lb_n)
						);
//M_MOD COUNTER		
mod_m_count device1(.clk(clk), .reset(rst_pulse), .count(), .pulse(pulse));  //m_mod counter set to 50ms delay = 54 minutes

always@(posedge clk, negedge reset_n)
begin
	if (!reset_n)
		begin
			state_reg = state_idle;
			count_reg = 0;
		end
	else
		begin
			state_reg <= state_next;
			count_reg <= count_next;
		end
end


//next state logic and outputs
always@*
begin
	start_n = 1'b1;
	rw = 1'b1;
	state_next = state_reg;
	count_next = count_reg;
	rst_pulse = 1'b1;
	case(state_reg)
	state_idle:
		begin
			if (write == 1'b0)
				begin
					state_next = state_write1;
					count_next = 0;
				end
			else
				if(read == 1'b0)
					begin
						state_next = state_read1;
						count_next = 0;
					end
		end //end state_idle	
	state_write1:
		begin
			rw = 1'b0;
			start_n = 1'b0;
			state_next = state_write2;
		end //end state_write1
	state_write2:
		begin
			rw = 1'b0;
			if (ready == 1)
				begin
				count_next = count_reg + 1'b1;
					if(count_next == 0)
						state_next = state_idle;
					else
						state_next = state_write1;
				end
			else
				state_next = state_write2;
		end //end state_write2
	state_read1:
		begin
			rw = 1'b1;
			start_n = 1'b0;
			state_next = state_read2;
			rst_pulse = 1'b0;
		end //end state_read1
	state_read2:
		begin
			rw = 1'b1;
			if ((ready == 1'b1) && (pulse == 1'b1))
				begin
				count_next = count_reg + 1'b1;
					if(count_next == 0)
						state_next = state_idle;
					else
						state_next = state_read1;
				end
			else
				state_next = state_read2;
		end //end state_read2
	default: state_next = state_reg;
   endcase
end

// data outputs
assign ledg = data_read[7:0];
assign ledr = data_read[15:8];  

endmodule

/*  SRAM CONTOLLER v2.0
**************************************************************** 
Summary:  a low level driver to fascillitate interaction
between an SRAM device and other peripherals.
*/

module sram_ctrl
(
//inputs
input wire clk , reset_n ,
input wire start_n, rw,
input wire [17:0] addr_in,
input wire [15:0] data_write,
//outputs
output reg ready,
output wire [15:0] data_read ,
output wire [17:0] sram_addr ,
output wire we_n, oe_n,
output wire ce_a_n , ub_a_n, lb_a_n,
//inout
inout wire [15:0] data_io
);

//states
localparam [1:0]  state_idle  = 3'b00,
						state_read  = 3'b01,
						state_write = 3'b10;
						
reg [2:0]   state_reg, state_next;
reg [15:0]  data_write_reg,   data_write_next;
reg [15:0]  data_read_reg, data_read_next;
reg [17:0]  addr_reg, addr_next;
reg we_next, oe_next, tri_next;
reg we_reg, oe_reg, tri_reg;

always@(posedge clk, negedge reset_n)
if(!reset_n)
	begin
		state_reg <= state_idle;
		addr_reg <= 0;
		data_write_reg <= 0;
		data_read_reg <= 0;
		we_reg <= 1'b1;
		oe_reg <= 1'b1;
		tri_reg <= 1'b1;
	end
else
	begin
		state_reg <= state_next;
		addr_reg  <= addr_next;
		data_write_reg <= data_write_next;
		data_read_reg <= data_read_next;
		we_reg <= we_next;
		oe_reg <= oe_next;
		tri_reg <= tri_next;
	end
		
//next state values and outputs
always@*
begin
	//default values
	addr_next = addr_reg;
	data_write_next = data_write_reg;
	data_read_next = data_read_reg;
	ready = 1'b0;
	oe_next = 1'b1;
	we_next = 1'b1;
	tri_next = 1'b1;
	//state machine
case(state_reg)		
	state_idle:
	begin
		ready = 1'b1;
		oe_next = 1'b1;
		if(start_n)  						
			state_next = state_reg;
		else
			begin
			  addr_next = addr_in;
			  if(rw == 1)
				begin
					state_next = state_read;  //BEGIN READ PROCESS
					oe_next = 1'b0;   
				end	
			  else
			   begin  								
					state_next = state_write;	// BEGIN WRITE PROCESS
					data_write_next = data_write;
					we_next = 1'b0;
					tri_next = 1'b0;
				end
			end
	end
	state_read:
		begin
			state_next = state_idle;
			data_read_next = data_io;
			oe_next = 1'b1;
		end
	state_write:
		begin
			state_next = state_idle;
			tri_next = 1'b0;
		end
	default: 
		state_next = state_idle;
endcase
end

//outputs
assign ce_a_n = 1'b0; 
assign ub_a_n = 1'b0;
assign lb_a_n = 1'b0;
assign oe_n = oe_reg;
assign we_n = we_reg;
assign sram_addr = addr_reg;
assign data_read = data_read_reg;

assign data_io =  (!tri_reg) ? data_write_reg : 16'bz;
endmodule


//*************************************************************************
//*************************************************************************
//*************************************************************************
//*************************************************************************
//*************************************************************************
module  mod_m_count
#(parameter M=50000) //2500000 = 50 ms | 250000 = 5 ms | 25000 = 500 us | 50000 = 1 ms
(
input  wire clk, reset,
output reg [log2(M)-1:0] count,
output wire pulse
);

localparam N = log2(M);
wire [N-1:0] count_next;

always@(posedge clk, negedge reset)
begin
	if(!reset)
		count <= 0;
	else 
		count <= count_next;
end

//next_state
assign count_next = (count == M-1) ? 0 : count + 1'b1;
//output
assign pulse = (count == M-1) ? 1'b1 : 1'b0;
//function
function integer log2(input integer m);
integer i;
begin
	log2 = 1;
	for (i=0; 2**i < m ;i=i+1)
		log2 = i + 1;
end
endfunction
endmodule
